module main;
  initial begin
    $display("С днем рождения. Желаю тебе  счастья, здоровья, успеха по жизни и в работе"); // non_trivial_congratulations
    $display("И пусть следующий тортик будет от Intel, вместе с предложением о сотрудничестве"); // dream_company
    $display("Уверен, у тебя все получится!");
  end
endmodule
